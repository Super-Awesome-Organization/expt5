// Group 2: Raj Patel, Zachary Rouviere, Evan Waxman
// Experiement 5 Part 1
// 9/24/21

// Description:
//	
`timescale 1ns/1ns

module  temp_to_led ( 
	input				clk,
	input				rst,
	output reg	[7:0]	led
);



        
endmodule
